library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

entity top_level_NCO_i2s_oscillator is 
port ( iReset : in std_logic := '0';
       iClock50Mhz : in std_logic := '0';
       oMasterClock : out std_logic := '0';
       oLeftRightClock : out std_logic := '0'; -- word select
       oSerialBitClock : out std_logic := '0'; -- sclk, bck. clock for data
       oData : out std_logic := '0'
       );
end entity;


architecture rtl of top_level_NCO_i2s_oscillator is
constant phaseInc : std_logic_vector (31 downto 0) := std_logic_vector(to_unsigned(85899,32)); -- 1000 Hz / 50000000Hz * 2^32
signal sSineNumber : std_logic_vector(15 downto 0);
signal mySignalL : std_logic_vector (23 downto 0) := (others => '0');
signal mySignalR : std_logic_vector (23 downto 0) := (others => '0');
signal sLeftRight : std_logic := '0';
begin
  waveform_generator : entity work.waveform_gen_14addr_16value(rtl)
  port map(clk => iClock50Mhz,
           reset => iReset,
	   sin_out => sSineNumber,
	   phase_inc => phaseInc);

   i2s_transmiter : entity work.i2s_master(rtl)
   generic map(CLK_FREQ => 50000000)
   port map(reset => not iReset,
            clk => iClock50Mhz,
	    mClk =>oMasterClock,
	    lrclk => sLeftRight,
	    sclk => oSerialBitClock,
	    sdata => oData,
	    data_l => mySignalL,
	    data_r => mySignalR);
   oLeftRightClock <= sLeftRight;
   mySignalL (23 downto 8) <= sSineNumber;
   mySignalR (23 downto 8) <= sSineNumber;
end rtl;
